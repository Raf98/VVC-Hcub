-- DST-VII 1D 8x8 utilizando MCU com Hcub para a multiplicação
-- e Macro Function para as somas
-- Rafael Santos; André Marcelo Coelho da Silva
-- Created: 18/12/2023


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


	
entity DST7_DCT8_32x32 is
	generic(
		Nbits				:  integer := 9;
		inBits			:  integer := 9;
		numInOutputs	:  integer := 64;
		outBits			:  integer := 19; --19 downto 0 -> 20 bits
		rNum				:  integer := 4;
		numTr				:  integer := 2
	);
	port(
		op:												 in std_logic;
		x0 ,x1 ,x2 ,x3 ,x4 ,x5 ,x6 ,x7: 			 in std_logic_vector(inBits - 1 downto 0);
		x8 ,x9 ,x10 ,x11 ,x12 ,x13 ,x14 ,x15:   in std_logic_vector(inBits - 1 downto 0);
		x16 ,x17 ,x18 ,x19 ,x20 ,x21 ,x22 ,x23: in std_logic_vector(inBits - 1 downto 0);
		x24 ,x25 ,x26 ,x27 ,x28 ,x29 ,x30 ,x31: in std_logic_vector(inBits - 1 downto 0);
		x32 ,x33 ,x34 ,x35 ,x36 ,x37 ,x38 ,x39: in std_logic_vector(inBits - 1 downto 0);
		x40 ,x41 ,x42 ,x43 ,x44 ,x45 ,x46 ,x47: in std_logic_vector(inBits - 1 downto 0);
		x48 ,x49 ,x50 ,x51 ,x52 ,x53 ,x54 ,x55: in std_logic_vector(inBits - 1 downto 0);
		x56 ,x57 ,x58 ,x59 ,x60 ,x61 ,x62 ,x63: in std_logic_vector(inBits - 1 downto 0);
		
		y0, y1, y2, y3, y4, y5, y6, y7		  : out std_logic_vector(outBits   downto 0);
		y8, y9, y10, y11, y12, y13, y14, y15  : out std_logic_vector(outBits   downto 0);
		y16, y17, y18, y19, y20, y21, y22, y23: out std_logic_vector(outBits   downto 0);
		y24, y25, y26, y27, y28, y29, y30, y31: out std_logic_vector(outBits   downto 0);
		y32, y33, y34, y35, y36, y37, y38, y39: out std_logic_vector(outBits   downto 0);
		y40, y41, y42, y43, y44, y45, y46, y47: out std_logic_vector(outBits   downto 0);
		y48, y49, y50, y51, y52, y53, y54, y55: out std_logic_vector(outBits   downto 0);
		y56, y57, y58, y59, y60, y61, y62, y63: out std_logic_vector(outBits   downto 0)
);

end DST7_DCT8_32x32;


architecture behavior of DST7_DCT8_32x32 is
		
		Component MCUHcub_DST7_DCT8_32x32 is
			PORT(
				x 		: in  std_logic_vector (inBits - 1  downto 0);
				x4  	: out std_logic_vector (outBits 	downto 0);
				x9  	: out std_logic_vector (outBits 	downto 0);
				x13 	: out std_logic_vector (outBits 	downto 0);
				x17 	: out std_logic_vector (outBits 	downto 0);
				x21 	: out std_logic_vector (outBits 	downto 0);
				x26 	: out std_logic_vector (outBits 	downto 0);
				x30 	: out std_logic_vector (outBits 	downto 0);
				x34 	: out std_logic_vector (outBits 	downto 0);
				x38 	: out std_logic_vector (outBits 	downto 0);
				x42 	: out std_logic_vector (outBits 	downto 0);
				x46 	: out std_logic_vector (outBits 	downto 0);
				x50 	: out std_logic_vector (outBits 	downto 0);
				x53 	: out std_logic_vector (outBits 	downto 0);
				x56 	: out std_logic_vector (outBits 	downto 0);
				x60 	: out std_logic_vector (outBits 	downto 0);
				x63 	: out std_logic_vector (outBits 	downto 0);
				x66 	: out std_logic_vector (outBits 	downto 0);
				x68 	: out std_logic_vector (outBits 	downto 0);
				x72 	: out std_logic_vector (outBits 	downto 0);
				x74 	: out std_logic_vector (outBits 	downto 0);
				x77 	: out std_logic_vector (outBits 	downto 0);
				x78 	: out std_logic_vector (outBits 	downto 0);
				x80 	: out std_logic_vector (outBits 	downto 0);
				x82 	: out std_logic_vector (outBits 	downto 0);
				x84 	: out std_logic_vector (outBits 	downto 0);
				x85 	: out std_logic_vector (outBits 	downto 0);
				x86 	: out std_logic_vector (outBits 	downto 0);
				x87 	: out std_logic_vector (outBits 	downto 0);
				x88 	: out std_logic_vector (outBits 	downto 0);
				x89 	: out std_logic_vector (outBits 	downto 0);
				x90 	: out std_logic_vector (outBits 	downto 0) 
			);
		end Component;
		
		
		type hcubOutputs is array( 0 to numInOutputs - 1 ) of std_logic_vector( outBits downto 0 );
		signal x_4, x_9, x_13, x_17, x_21, x_26, x_30, x_34, x_38, x_42, x_46, x_50, x_53, x_56, x_60, x_63: hcubOutputs;
		signal x_66, x_68, x_72, x_74, x_77, x_78, x_80, x_82, x_84, x_85, x_86, x_87, x_88, x_89, x_90		: hcubOutputs;
		
		type inputSignals is array( 0 to numInOutputs - 1 ) of std_logic_vector( inBits - 1 downto 0 );
		signal x: inputSignals;
		
		type outputSignals is array( 0 to numInOutputs - 1 ) of std_logic_vector( outBits downto 0 );
		signal y, y_dct, y_dst: outputSignals;
	

begin 
x(0) <= x0;
x(1) <= x1;
x(2) <= x2;
x(3) <= x3;
x(4) <= x4;
x(5) <= x5;
x(6) <= x6;
x(7) <= x7;
x(8) <= x8;
x(9) <= x9;
x(10) <= x10;
x(11) <= x11;
x(12) <= x12;
x(13) <= x13;
x(14) <= x14;
x(15) <= x15;
x(16) <= x16;
x(17) <= x17;
x(18) <= x18;
x(19) <= x19;
x(20) <= x20;
x(21) <= x21;
x(22) <= x22;
x(23) <= x23;
x(24) <= x24;
x(25) <= x25;
x(26) <= x26;
x(27) <= x27;
x(28) <= x28;
x(29) <= x29;
x(30) <= x30;
x(31) <= x31;
x(32) <= x32;
x(33) <= x33;
x(34) <= x34;
x(35) <= x35;
x(36) <= x36;
x(37) <= x37;
x(38) <= x38;
x(39) <= x39;
x(40) <= x40;
x(41) <= x41;
x(42) <= x42;
x(43) <= x43;
x(44) <= x44;
x(45) <= x45;
x(46) <= x46;
x(47) <= x47;
x(48) <= x48;
x(49) <= x49;
x(50) <= x50;
x(51) <= x51;
x(52) <= x52;
x(53) <= x53;
x(54) <= x54;
x(55) <= x55;
x(56) <= x56;
x(57) <= x57;
x(58) <= x58;
x(59) <= x59;
x(60) <= x60;
x(61) <= x61;
x(62) <= x62;
x(63) <= x63;


			generateMCUs:        
            for i in 0 to numInOutputs-1 generate
						  
					MCU: MCUHcub_DST7_DCT8_32x32 
					port map(
						x 	 => x(i),
						x4  => x_4(i),
						x9  => x_9(i),
						x13 => x_13(i),
						x17 => x_17(i),
						x21 => x_21(i),
						x26 => x_26(i),
						x30 => x_30(i),
						x34 => x_34(i),
						x38 => x_38(i),
						x42 => x_42(i),
						x46 => x_46(i),
						x50 => x_50(i),
						x53 => x_53(i),
						x56 => x_56(i),
						x60 => x_60(i),
						x63 => x_63(i),
						x66 => x_66(i),
						x68 => x_68(i),
						x72 => x_72(i),
						x74 => x_74(i),
						x77 => x_77(i),
						x78 => x_78(i),
						x80 => x_80(i),
						x82 => x_82(i),
						x84 => x_84(i),
						x85 => x_85(i),
						x86 => x_86(i),
						x87 => x_87(i),
						x88 => x_88(i),
						x89 => x_89(i),
						x90 => x_90(i));
						  
				end generate generateMCUs;
        
        generateSignalsOutputsDCT8:        
            for i in 0 to numTr - 1 generate

						y_dct(i*32 + 0) <= x_90(i*32 + 0) + x_90(i*32 + 1) + x_89(i*32 + 2) + x_88(i*32 + 3) + x_87(i*32 + 4) + x_86(i*32 + 5) + x_85(i*32 + 6) + x_84(i*32 + 7) + x_82(i*32 + 8) + x_80(i*32 + 9) + x_78(i*32 + 10) + x_77(i*32 + 11) + x_74(i*32 + 12) + x_72(i*32 + 13) + x_68(i*32 + 14) + x_66(i*32 + 15) + x_63(i*32 + 16) + x_60(i*32 + 17) + x_56(i*32 + 18) + x_53(i*32 + 19) + x_50(i*32 + 20) + x_46(i*32 + 21) + x_42(i*32 + 22) + x_38(i*32 + 23) + x_34(i*32 + 24) + x_30(i*32 + 25) + x_26(i*32 + 26) + x_21(i*32 + 27) + x_17(i*32 + 28) + x_13(i*32 + 29) + x_9(i*32 + 30) + x_4(i*32 + 31);
						y_dct(i*32 + 1) <= x_90(i*32 + 0) + x_87(i*32 + 1) + x_84(i*32 + 2) + x_78(i*32 + 3) + x_72(i*32 + 4) + x_63(i*32 + 5) + x_53(i*32 + 6) + x_42(i*32 + 7) + x_30(i*32 + 8) + x_17(i*32 + 9) + x_4(i*32 + 10) - x_9(i*32 + 11) - x_21(i*32 + 12) - x_34(i*32 + 13) - x_46(i*32 + 14) - x_56(i*32 + 15) - x_66(i*32 + 16) - x_74(i*32 + 17) - x_80(i*32 + 18) - x_85(i*32 + 19) - x_88(i*32 + 20) - x_90(i*32 + 21) - x_89(i*32 + 22) - x_86(i*32 + 23) - x_82(i*32 + 24) - x_77(i*32 + 25) - x_68(i*32 + 26) - x_60(i*32 + 27) - x_50(i*32 + 28) - x_38(i*32 + 29) - x_26(i*32 + 30) - x_13(i*32 + 31);
						y_dct(i*32 + 2) <= x_89(i*32 + 0) + x_84(i*32 + 1) + x_74(i*32 + 2) + x_60(i*32 + 3) + x_42(i*32 + 4) + x_21(i*32 + 5) - x_21(i*32 + 7) - x_42(i*32 + 8) - x_60(i*32 + 9) - x_74(i*32 + 10) - x_84(i*32 + 11) - x_89(i*32 + 12) - x_89(i*32 + 13) - x_84(i*32 + 14) - x_74(i*32 + 15) - x_60(i*32 + 16) - x_42(i*32 + 17) - x_21(i*32 + 18) + x_21(i*32 + 20) + x_42(i*32 + 21) + x_60(i*32 + 22) + x_74(i*32 + 23) + x_84(i*32 + 24) + x_89(i*32 + 25) + x_89(i*32 + 26) + x_84(i*32 + 27) + x_74(i*32 + 28) + x_60(i*32 + 29) + x_42(i*32 + 30) + x_21(i*32 + 31);
						y_dct(i*32 + 3) <= x_88(i*32 + 0) + x_78(i*32 + 1) + x_60(i*32 + 2) + x_34(i*32 + 3) + x_4(i*32 + 4) - x_26(i*32 + 5) - x_53(i*32 + 6) - x_74(i*32 + 7) - x_86(i*32 + 8) - x_90(i*32 + 9) - x_82(i*32 + 10) - x_66(i*32 + 11) - x_42(i*32 + 12) - x_13(i*32 + 13) + x_17(i*32 + 14) + x_46(i*32 + 15) + x_68(i*32 + 16) + x_84(i*32 + 17) + x_90(i*32 + 18) + x_85(i*32 + 19) + x_72(i*32 + 20) + x_50(i*32 + 21) + x_21(i*32 + 22) - x_9(i*32 + 23) - x_38(i*32 + 24) - x_63(i*32 + 25) - x_80(i*32 + 26) - x_89(i*32 + 27) - x_87(i*32 + 28) - x_77(i*32 + 29) - x_56(i*32 + 30) - x_30(i*32 + 31);
						y_dct(i*32 + 4) <= x_87(i*32 + 0) + x_72(i*32 + 1) + x_42(i*32 + 2) + x_4(i*32 + 3) - x_34(i*32 + 4) - x_66(i*32 + 5) - x_85(i*32 + 6) - x_89(i*32 + 7) - x_77(i*32 + 8) - x_50(i*32 + 9) - x_13(i*32 + 10) + x_26(i*32 + 11) + x_60(i*32 + 12) + x_82(i*32 + 13) + x_90(i*32 + 14) + x_80(i*32 + 15) + x_56(i*32 + 16) + x_21(i*32 + 17) - x_17(i*32 + 18) - x_53(i*32 + 19) - x_78(i*32 + 20) - x_90(i*32 + 21) - x_84(i*32 + 22) - x_63(i*32 + 23) - x_30(i*32 + 24) + x_9(i*32 + 25) + x_46(i*32 + 26) + x_74(i*32 + 27) + x_88(i*32 + 28) + x_86(i*32 + 29) + x_68(i*32 + 30) + x_38(i*32 + 31);
						y_dct(i*32 + 5) <= x_86(i*32 + 0) + x_63(i*32 + 1) + x_21(i*32 + 2) - x_26(i*32 + 3) - x_66(i*32 + 4) - x_87(i*32 + 5) - x_85(i*32 + 6) - x_60(i*32 + 7) - x_17(i*32 + 8) + x_30(i*32 + 9) + x_68(i*32 + 10) + x_88(i*32 + 11) + x_84(i*32 + 12) + x_56(i*32 + 13) + x_13(i*32 + 14) - x_34(i*32 + 15) - x_72(i*32 + 16) - x_89(i*32 + 17) - x_82(i*32 + 18) - x_53(i*32 + 19) - x_9(i*32 + 20) + x_38(i*32 + 21) + x_74(i*32 + 22) + x_90(i*32 + 23) + x_80(i*32 + 24) + x_50(i*32 + 25) + x_4(i*32 + 26) - x_42(i*32 + 27) - x_77(i*32 + 28) - x_90(i*32 + 29) - x_78(i*32 + 30) - x_46(i*32 + 31);
						y_dct(i*32 + 6) <= x_85(i*32 + 0) + x_53(i*32 + 1) - x_53(i*32 + 3) - x_85(i*32 + 4) - x_85(i*32 + 5) - x_53(i*32 + 6) + x_53(i*32 + 8) + x_85(i*32 + 9) + x_85(i*32 + 10) + x_53(i*32 + 11) - x_53(i*32 + 13) - x_85(i*32 + 14) - x_85(i*32 + 15) - x_53(i*32 + 16) + x_53(i*32 + 18) + x_85(i*32 + 19) + x_85(i*32 + 20) + x_53(i*32 + 21) - x_53(i*32 + 23) - x_85(i*32 + 24) - x_85(i*32 + 25) - x_53(i*32 + 26) + x_53(i*32 + 28) + x_85(i*32 + 29) + x_85(i*32 + 30) + x_53(i*32 + 31);
						y_dct(i*32 + 7) <= x_84(i*32 + 0) + x_42(i*32 + 1) - x_21(i*32 + 2) - x_74(i*32 + 3) - x_89(i*32 + 4) - x_60(i*32 + 5) + x_60(i*32 + 7) + x_89(i*32 + 8) + x_74(i*32 + 9) + x_21(i*32 + 10) - x_42(i*32 + 11) - x_84(i*32 + 12) - x_84(i*32 + 13) - x_42(i*32 + 14) + x_21(i*32 + 15) + x_74(i*32 + 16) + x_89(i*32 + 17) + x_60(i*32 + 18) - x_60(i*32 + 20) - x_89(i*32 + 21) - x_74(i*32 + 22) - x_21(i*32 + 23) + x_42(i*32 + 24) + x_84(i*32 + 25) + x_84(i*32 + 26) + x_42(i*32 + 27) - x_21(i*32 + 28) - x_74(i*32 + 29) - x_89(i*32 + 30) - x_60(i*32 + 31);
						y_dct(i*32 + 8) <= x_82(i*32 + 0) + x_30(i*32 + 1) - x_42(i*32 + 2) - x_86(i*32 + 3) - x_77(i*32 + 4) - x_17(i*32 + 5) + x_53(i*32 + 6) + x_89(i*32 + 7) + x_68(i*32 + 8) + x_4(i*32 + 9) - x_63(i*32 + 10) - x_90(i*32 + 11) - x_60(i*32 + 12) + x_9(i*32 + 13) + x_72(i*32 + 14) + x_88(i*32 + 15) + x_50(i*32 + 16) - x_21(i*32 + 17) - x_78(i*32 + 18) - x_85(i*32 + 19) - x_38(i*32 + 20) + x_34(i*32 + 21) + x_84(i*32 + 22) + x_80(i*32 + 23) + x_26(i*32 + 24) - x_46(i*32 + 25) - x_87(i*32 + 26) - x_74(i*32 + 27) - x_13(i*32 + 28) + x_56(i*32 + 29) + x_90(i*32 + 30) + x_66(i*32 + 31);
						y_dct(i*32 + 9) <= x_80(i*32 + 0) + x_17(i*32 + 1) - x_60(i*32 + 2) - x_90(i*32 + 3) - x_50(i*32 + 4) + x_30(i*32 + 5) + x_85(i*32 + 6) + x_74(i*32 + 7) + x_4(i*32 + 8) - x_68(i*32 + 9) - x_87(i*32 + 10) - x_38(i*32 + 11) + x_42(i*32 + 12) + x_88(i*32 + 13) + x_66(i*32 + 14) - x_9(i*32 + 15) - x_77(i*32 + 16) - x_84(i*32 + 17) - x_26(i*32 + 18) + x_53(i*32 + 19) + x_90(i*32 + 20) + x_56(i*32 + 21) - x_21(i*32 + 22) - x_82(i*32 + 23) - x_78(i*32 + 24) - x_13(i*32 + 25) + x_63(i*32 + 26) + x_89(i*32 + 27) + x_46(i*32 + 28) - x_34(i*32 + 29) - x_86(i*32 + 30) - x_72(i*32 + 31);
						y_dct(i*32 + 10) <= x_78(i*32 + 0) + x_4(i*32 + 1) - x_74(i*32 + 2) - x_82(i*32 + 3) - x_13(i*32 + 4) + x_68(i*32 + 5) + x_85(i*32 + 6) + x_21(i*32 + 7) - x_63(i*32 + 8) - x_87(i*32 + 9) - x_30(i*32 + 10) + x_56(i*32 + 11) + x_89(i*32 + 12) + x_38(i*32 + 13) - x_50(i*32 + 14) - x_90(i*32 + 15) - x_46(i*32 + 16) + x_42(i*32 + 17) + x_90(i*32 + 18) + x_53(i*32 + 19) - x_34(i*32 + 20) - x_88(i*32 + 21) - x_60(i*32 + 22) + x_26(i*32 + 23) + x_86(i*32 + 24) + x_66(i*32 + 25) - x_17(i*32 + 26) - x_84(i*32 + 27) - x_72(i*32 + 28) + x_9(i*32 + 29) + x_80(i*32 + 30) + x_77(i*32 + 31);
						y_dct(i*32 + 11) <= x_77(i*32 + 0) - x_9(i*32 + 1) - x_84(i*32 + 2) - x_66(i*32 + 3) + x_26(i*32 + 4) + x_88(i*32 + 5) + x_53(i*32 + 6) - x_42(i*32 + 7) - x_90(i*32 + 8) - x_38(i*32 + 9) + x_56(i*32 + 10) + x_87(i*32 + 11) + x_21(i*32 + 12) - x_68(i*32 + 13) - x_82(i*32 + 14) - x_4(i*32 + 15) + x_78(i*32 + 16) + x_74(i*32 + 17) - x_13(i*32 + 18) - x_85(i*32 + 19) - x_63(i*32 + 20) + x_30(i*32 + 21) + x_89(i*32 + 22) + x_50(i*32 + 23) - x_46(i*32 + 24) - x_90(i*32 + 25) - x_34(i*32 + 26) + x_60(i*32 + 27) + x_86(i*32 + 28) + x_17(i*32 + 29) - x_72(i*32 + 30) - x_80(i*32 + 31);
						y_dct(i*32 + 12) <= x_74(i*32 + 0) - x_21(i*32 + 1) - x_89(i*32 + 2) - x_42(i*32 + 3) + x_60(i*32 + 4) + x_84(i*32 + 5) - x_84(i*32 + 7) - x_60(i*32 + 8) + x_42(i*32 + 9) + x_89(i*32 + 10) + x_21(i*32 + 11) - x_74(i*32 + 12) - x_74(i*32 + 13) + x_21(i*32 + 14) + x_89(i*32 + 15) + x_42(i*32 + 16) - x_60(i*32 + 17) - x_84(i*32 + 18) + x_84(i*32 + 20) + x_60(i*32 + 21) - x_42(i*32 + 22) - x_89(i*32 + 23) - x_21(i*32 + 24) + x_74(i*32 + 25) + x_74(i*32 + 26) - x_21(i*32 + 27) - x_89(i*32 + 28) - x_42(i*32 + 29) + x_60(i*32 + 30) + x_84(i*32 + 31);
						y_dct(i*32 + 13) <= x_72(i*32 + 0) - x_34(i*32 + 1) - x_89(i*32 + 2) - x_13(i*32 + 3) + x_82(i*32 + 4) + x_56(i*32 + 5) - x_53(i*32 + 6) - x_84(i*32 + 7) + x_9(i*32 + 8) + x_88(i*32 + 9) + x_38(i*32 + 10) - x_68(i*32 + 11) - x_74(i*32 + 12) + x_30(i*32 + 13) + x_90(i*32 + 14) + x_17(i*32 + 15) - x_80(i*32 + 16) - x_60(i*32 + 17) + x_50(i*32 + 18) + x_85(i*32 + 19) - x_4(i*32 + 20) - x_87(i*32 + 21) - x_42(i*32 + 22) + x_66(i*32 + 23) + x_77(i*32 + 24) - x_26(i*32 + 25) - x_90(i*32 + 26) - x_21(i*32 + 27) + x_78(i*32 + 28) + x_63(i*32 + 29) - x_46(i*32 + 30) - x_86(i*32 + 31);
						y_dct(i*32 + 14) <= x_68(i*32 + 0) - x_46(i*32 + 1) - x_84(i*32 + 2) + x_17(i*32 + 3) + x_90(i*32 + 4) + x_13(i*32 + 5) - x_85(i*32 + 6) - x_42(i*32 + 7) + x_72(i*32 + 8) + x_66(i*32 + 9) - x_50(i*32 + 10) - x_82(i*32 + 11) + x_21(i*32 + 12) + x_90(i*32 + 13) + x_9(i*32 + 14) - x_86(i*32 + 15) - x_38(i*32 + 16) + x_74(i*32 + 17) + x_63(i*32 + 18) - x_53(i*32 + 19) - x_80(i*32 + 20) + x_26(i*32 + 21) + x_89(i*32 + 22) + x_4(i*32 + 23) - x_87(i*32 + 24) - x_34(i*32 + 25) + x_77(i*32 + 26) + x_60(i*32 + 27) - x_56(i*32 + 28) - x_78(i*32 + 29) + x_30(i*32 + 30) + x_88(i*32 + 31);
						y_dct(i*32 + 15) <= x_66(i*32 + 0) - x_56(i*32 + 1) - x_74(i*32 + 2) + x_46(i*32 + 3) + x_80(i*32 + 4) - x_34(i*32 + 5) - x_85(i*32 + 6) + x_21(i*32 + 7) + x_88(i*32 + 8) - x_9(i*32 + 9) - x_90(i*32 + 10) - x_4(i*32 + 11) + x_89(i*32 + 12) + x_17(i*32 + 13) - x_86(i*32 + 14) - x_30(i*32 + 15) + x_82(i*32 + 16) + x_42(i*32 + 17) - x_77(i*32 + 18) - x_53(i*32 + 19) + x_68(i*32 + 20) + x_63(i*32 + 21) - x_60(i*32 + 22) - x_72(i*32 + 23) + x_50(i*32 + 24) + x_78(i*32 + 25) - x_38(i*32 + 26) - x_84(i*32 + 27) + x_26(i*32 + 28) + x_87(i*32 + 29) - x_13(i*32 + 30) - x_90(i*32 + 31);
						y_dct(i*32 + 16) <= x_63(i*32 + 0) - x_66(i*32 + 1) - x_60(i*32 + 2) + x_68(i*32 + 3) + x_56(i*32 + 4) - x_72(i*32 + 5) - x_53(i*32 + 6) + x_74(i*32 + 7) + x_50(i*32 + 8) - x_77(i*32 + 9) - x_46(i*32 + 10) + x_78(i*32 + 11) + x_42(i*32 + 12) - x_80(i*32 + 13) - x_38(i*32 + 14) + x_82(i*32 + 15) + x_34(i*32 + 16) - x_84(i*32 + 17) - x_30(i*32 + 18) + x_85(i*32 + 19) + x_26(i*32 + 20) - x_86(i*32 + 21) - x_21(i*32 + 22) + x_87(i*32 + 23) + x_17(i*32 + 24) - x_88(i*32 + 25) - x_13(i*32 + 26) + x_89(i*32 + 27) + x_9(i*32 + 28) - x_90(i*32 + 29) - x_4(i*32 + 30) + x_90(i*32 + 31);
						y_dct(i*32 + 17) <= x_60(i*32 + 0) - x_74(i*32 + 1) - x_42(i*32 + 2) + x_84(i*32 + 3) + x_21(i*32 + 4) - x_89(i*32 + 5) + x_89(i*32 + 7) - x_21(i*32 + 8) - x_84(i*32 + 9) + x_42(i*32 + 10) + x_74(i*32 + 11) - x_60(i*32 + 12) - x_60(i*32 + 13) + x_74(i*32 + 14) + x_42(i*32 + 15) - x_84(i*32 + 16) - x_21(i*32 + 17) + x_89(i*32 + 18) - x_89(i*32 + 20) + x_21(i*32 + 21) + x_84(i*32 + 22) - x_42(i*32 + 23) - x_74(i*32 + 24) + x_60(i*32 + 25) + x_60(i*32 + 26) - x_74(i*32 + 27) - x_42(i*32 + 28) + x_84(i*32 + 29) + x_21(i*32 + 30) - x_89(i*32 + 31);
						y_dct(i*32 + 18) <= x_56(i*32 + 0) - x_80(i*32 + 1) - x_21(i*32 + 2) + x_90(i*32 + 3) - x_17(i*32 + 4) - x_82(i*32 + 5) + x_53(i*32 + 6) + x_60(i*32 + 7) - x_78(i*32 + 8) - x_26(i*32 + 9) + x_90(i*32 + 10) - x_13(i*32 + 11) - x_84(i*32 + 12) + x_50(i*32 + 13) + x_63(i*32 + 14) - x_77(i*32 + 15) - x_30(i*32 + 16) + x_89(i*32 + 17) - x_9(i*32 + 18) - x_85(i*32 + 19) + x_46(i*32 + 20) + x_66(i*32 + 21) - x_74(i*32 + 22) - x_34(i*32 + 23) + x_88(i*32 + 24) - x_4(i*32 + 25) - x_86(i*32 + 26) + x_42(i*32 + 27) + x_68(i*32 + 28) - x_72(i*32 + 29) - x_38(i*32 + 30) + x_87(i*32 + 31);
						y_dct(i*32 + 19) <= x_53(i*32 + 0) - x_85(i*32 + 1) + x_85(i*32 + 3) - x_53(i*32 + 4) - x_53(i*32 + 5) + x_85(i*32 + 6) - x_85(i*32 + 8) + x_53(i*32 + 9) + x_53(i*32 + 10) - x_85(i*32 + 11) + x_85(i*32 + 13) - x_53(i*32 + 14) - x_53(i*32 + 15) + x_85(i*32 + 16) - x_85(i*32 + 18) + x_53(i*32 + 19) + x_53(i*32 + 20) - x_85(i*32 + 21) + x_85(i*32 + 23) - x_53(i*32 + 24) - x_53(i*32 + 25) + x_85(i*32 + 26) - x_85(i*32 + 28) + x_53(i*32 + 29) + x_53(i*32 + 30) - x_85(i*32 + 31);
						y_dct(i*32 + 20) <= x_50(i*32 + 0) - x_88(i*32 + 1) + x_21(i*32 + 2) + x_72(i*32 + 3) - x_78(i*32 + 4) - x_9(i*32 + 5) + x_85(i*32 + 6) - x_60(i*32 + 7) - x_38(i*32 + 8) + x_90(i*32 + 9) - x_34(i*32 + 10) - x_63(i*32 + 11) + x_84(i*32 + 12) - x_4(i*32 + 13) - x_80(i*32 + 14) + x_68(i*32 + 15) + x_26(i*32 + 16) - x_89(i*32 + 17) + x_46(i*32 + 18) + x_53(i*32 + 19) - x_87(i*32 + 20) + x_17(i*32 + 21) + x_74(i*32 + 22) - x_77(i*32 + 23) - x_13(i*32 + 24) + x_86(i*32 + 25) - x_56(i*32 + 26) - x_42(i*32 + 27) + x_90(i*32 + 28) - x_30(i*32 + 29) - x_66(i*32 + 30) + x_82(i*32 + 31);
						y_dct(i*32 + 21) <= x_46(i*32 + 0) - x_90(i*32 + 1) + x_42(i*32 + 2) + x_50(i*32 + 3) - x_90(i*32 + 4) + x_38(i*32 + 5) + x_53(i*32 + 6) - x_89(i*32 + 7) + x_34(i*32 + 8) + x_56(i*32 + 9) - x_88(i*32 + 10) + x_30(i*32 + 11) + x_60(i*32 + 12) - x_87(i*32 + 13) + x_26(i*32 + 14) + x_63(i*32 + 15) - x_86(i*32 + 16) + x_21(i*32 + 17) + x_66(i*32 + 18) - x_85(i*32 + 19) + x_17(i*32 + 20) + x_68(i*32 + 21) - x_84(i*32 + 22) + x_13(i*32 + 23) + x_72(i*32 + 24) - x_82(i*32 + 25) + x_9(i*32 + 26) + x_74(i*32 + 27) - x_80(i*32 + 28) + x_4(i*32 + 29) + x_77(i*32 + 30) - x_78(i*32 + 31);
						y_dct(i*32 + 22) <= x_42(i*32 + 0) - x_89(i*32 + 1) + x_60(i*32 + 2) + x_21(i*32 + 3) - x_84(i*32 + 4) + x_74(i*32 + 5) - x_74(i*32 + 7) + x_84(i*32 + 8) - x_21(i*32 + 9) - x_60(i*32 + 10) + x_89(i*32 + 11) - x_42(i*32 + 12) - x_42(i*32 + 13) + x_89(i*32 + 14) - x_60(i*32 + 15) - x_21(i*32 + 16) + x_84(i*32 + 17) - x_74(i*32 + 18) + x_74(i*32 + 20) - x_84(i*32 + 21) + x_21(i*32 + 22) + x_60(i*32 + 23) - x_89(i*32 + 24) + x_42(i*32 + 25) + x_42(i*32 + 26) - x_89(i*32 + 27) + x_60(i*32 + 28) + x_21(i*32 + 29) - x_84(i*32 + 30) + x_74(i*32 + 31);
						y_dct(i*32 + 23) <= x_38(i*32 + 0) - x_86(i*32 + 1) + x_74(i*32 + 2) - x_9(i*32 + 3) - x_63(i*32 + 4) + x_90(i*32 + 5) - x_53(i*32 + 6) - x_21(i*32 + 7) + x_80(i*32 + 8) - x_82(i*32 + 9) + x_26(i*32 + 10) + x_50(i*32 + 11) - x_89(i*32 + 12) + x_66(i*32 + 13) + x_4(i*32 + 14) - x_72(i*32 + 15) + x_87(i*32 + 16) - x_42(i*32 + 17) - x_34(i*32 + 18) + x_85(i*32 + 19) - x_77(i*32 + 20) + x_13(i*32 + 21) + x_60(i*32 + 22) - x_90(i*32 + 23) + x_56(i*32 + 24) + x_17(i*32 + 25) - x_78(i*32 + 26) + x_84(i*32 + 27) - x_30(i*32 + 28) - x_46(i*32 + 29) + x_88(i*32 + 30) - x_68(i*32 + 31);
						y_dct(i*32 + 24) <= x_34(i*32 + 0) - x_82(i*32 + 1) + x_84(i*32 + 2) - x_38(i*32 + 3) - x_30(i*32 + 4) + x_80(i*32 + 5) - x_85(i*32 + 6) + x_42(i*32 + 7) + x_26(i*32 + 8) - x_78(i*32 + 9) + x_86(i*32 + 10) - x_46(i*32 + 11) - x_21(i*32 + 12) + x_77(i*32 + 13) - x_87(i*32 + 14) + x_50(i*32 + 15) + x_17(i*32 + 16) - x_74(i*32 + 17) + x_88(i*32 + 18) - x_53(i*32 + 19) - x_13(i*32 + 20) + x_72(i*32 + 21) - x_89(i*32 + 22) + x_56(i*32 + 23) + x_9(i*32 + 24) - x_68(i*32 + 25) + x_90(i*32 + 26) - x_60(i*32 + 27) - x_4(i*32 + 28) + x_66(i*32 + 29) - x_90(i*32 + 30) + x_63(i*32 + 31);
						y_dct(i*32 + 25) <= x_30(i*32 + 0) - x_77(i*32 + 1) + x_89(i*32 + 2) - x_63(i*32 + 3) + x_9(i*32 + 4) + x_50(i*32 + 5) - x_85(i*32 + 6) + x_84(i*32 + 7) - x_46(i*32 + 8) - x_13(i*32 + 9) + x_66(i*32 + 10) - x_90(i*32 + 11) + x_74(i*32 + 12) - x_26(i*32 + 13) - x_34(i*32 + 14) + x_78(i*32 + 15) - x_88(i*32 + 16) + x_60(i*32 + 17) - x_4(i*32 + 18) - x_53(i*32 + 19) + x_86(i*32 + 20) - x_82(i*32 + 21) + x_42(i*32 + 22) + x_17(i*32 + 23) - x_68(i*32 + 24) + x_90(i*32 + 25) - x_72(i*32 + 26) + x_21(i*32 + 27) + x_38(i*32 + 28) - x_80(i*32 + 29) + x_87(i*32 + 30) - x_56(i*32 + 31);
						y_dct(i*32 + 26) <= x_26(i*32 + 0) - x_68(i*32 + 1) + x_89(i*32 + 2) - x_80(i*32 + 3) + x_46(i*32 + 4) + x_4(i*32 + 5) - x_53(i*32 + 6) + x_84(i*32 + 7) - x_87(i*32 + 8) + x_63(i*32 + 9) - x_17(i*32 + 10) - x_34(i*32 + 11) + x_74(i*32 + 12) - x_90(i*32 + 13) + x_77(i*32 + 14) - x_38(i*32 + 15) - x_13(i*32 + 16) + x_60(i*32 + 17) - x_86(i*32 + 18) + x_85(i*32 + 19) - x_56(i*32 + 20) + x_9(i*32 + 21) + x_42(i*32 + 22) - x_78(i*32 + 23) + x_90(i*32 + 24) - x_72(i*32 + 25) + x_30(i*32 + 26) + x_21(i*32 + 27) - x_66(i*32 + 28) + x_88(i*32 + 29) - x_82(i*32 + 30) + x_50(i*32 + 31);
						y_dct(i*32 + 27) <= x_21(i*32 + 0) - x_60(i*32 + 1) + x_84(i*32 + 2) - x_89(i*32 + 3) + x_74(i*32 + 4) - x_42(i*32 + 5) + x_42(i*32 + 7) - x_74(i*32 + 8) + x_89(i*32 + 9) - x_84(i*32 + 10) + x_60(i*32 + 11) - x_21(i*32 + 12) - x_21(i*32 + 13) + x_60(i*32 + 14) - x_84(i*32 + 15) + x_89(i*32 + 16) - x_74(i*32 + 17) + x_42(i*32 + 18) - x_42(i*32 + 20) + x_74(i*32 + 21) - x_89(i*32 + 22) + x_84(i*32 + 23) - x_60(i*32 + 24) + x_21(i*32 + 25) + x_21(i*32 + 26) - x_60(i*32 + 27) + x_84(i*32 + 28) - x_89(i*32 + 29) + x_74(i*32 + 30) - x_42(i*32 + 31);
						y_dct(i*32 + 28) <= x_17(i*32 + 0) - x_50(i*32 + 1) + x_74(i*32 + 2) - x_87(i*32 + 3) + x_88(i*32 + 4) - x_77(i*32 + 5) + x_53(i*32 + 6) - x_21(i*32 + 7) - x_13(i*32 + 8) + x_46(i*32 + 9) - x_72(i*32 + 10) + x_86(i*32 + 11) - x_89(i*32 + 12) + x_78(i*32 + 13) - x_56(i*32 + 14) + x_26(i*32 + 15) + x_9(i*32 + 16) - x_42(i*32 + 17) + x_68(i*32 + 18) - x_85(i*32 + 19) + x_90(i*32 + 20) - x_80(i*32 + 21) + x_60(i*32 + 22) - x_30(i*32 + 23) - x_4(i*32 + 24) + x_38(i*32 + 25) - x_66(i*32 + 26) + x_84(i*32 + 27) - x_90(i*32 + 28) + x_82(i*32 + 29) - x_63(i*32 + 30) + x_34(i*32 + 31);
						y_dct(i*32 + 29) <= x_13(i*32 + 0) - x_38(i*32 + 1) + x_60(i*32 + 2) - x_77(i*32 + 3) + x_86(i*32 + 4) - x_90(i*32 + 5) + x_85(i*32 + 6) - x_74(i*32 + 7) + x_56(i*32 + 8) - x_34(i*32 + 9) + x_9(i*32 + 10) + x_17(i*32 + 11) - x_42(i*32 + 12) + x_63(i*32 + 13) - x_78(i*32 + 14) + x_87(i*32 + 15) - x_90(i*32 + 16) + x_84(i*32 + 17) - x_72(i*32 + 18) + x_53(i*32 + 19) - x_30(i*32 + 20) + x_4(i*32 + 21) + x_21(i*32 + 22) - x_46(i*32 + 23) + x_66(i*32 + 24) - x_80(i*32 + 25) + x_88(i*32 + 26) - x_89(i*32 + 27) + x_82(i*32 + 28) - x_68(i*32 + 29) + x_50(i*32 + 30) - x_26(i*32 + 31);
						y_dct(i*32 + 30) <= x_9(i*32 + 0) - x_26(i*32 + 1) + x_42(i*32 + 2) - x_56(i*32 + 3) + x_68(i*32 + 4) - x_78(i*32 + 5) + x_85(i*32 + 6) - x_89(i*32 + 7) + x_90(i*32 + 8) - x_86(i*32 + 9) + x_80(i*32 + 10) - x_72(i*32 + 11) + x_60(i*32 + 12) - x_46(i*32 + 13) + x_30(i*32 + 14) - x_13(i*32 + 15) - x_4(i*32 + 16) + x_21(i*32 + 17) - x_38(i*32 + 18) + x_53(i*32 + 19) - x_66(i*32 + 20) + x_77(i*32 + 21) - x_84(i*32 + 22) + x_88(i*32 + 23) - x_90(i*32 + 24) + x_87(i*32 + 25) - x_82(i*32 + 26) + x_74(i*32 + 27) - x_63(i*32 + 28) + x_50(i*32 + 29) - x_34(i*32 + 30) + x_17(i*32 + 31);
						y_dct(i*32 + 31) <= x_4(i*32 + 0) - x_13(i*32 + 1) + x_21(i*32 + 2) - x_30(i*32 + 3) + x_38(i*32 + 4) - x_46(i*32 + 5) + x_53(i*32 + 6) - x_60(i*32 + 7) + x_66(i*32 + 8) - x_72(i*32 + 9) + x_77(i*32 + 10) - x_80(i*32 + 11) + x_84(i*32 + 12) - x_86(i*32 + 13) + x_88(i*32 + 14) - x_90(i*32 + 15) + x_90(i*32 + 16) - x_89(i*32 + 17) + x_87(i*32 + 18) - x_85(i*32 + 19) + x_82(i*32 + 20) - x_78(i*32 + 21) + x_74(i*32 + 22) - x_68(i*32 + 23) + x_63(i*32 + 24) - x_56(i*32 + 25) + x_50(i*32 + 26) - x_42(i*32 + 27) + x_34(i*32 + 28) - x_26(i*32 + 29) + x_17(i*32 + 30) - x_9(i*32 + 31);
	  
            end generate generateSignalsOutputsDCT8;
				
				generateSignalsOutputsDST7:        
            for i in 0 to numTr - 1 generate
						
						y_dst(i*32 + 0) <= x_4(i*32 + 0) + x_13(i*32 + 1) + x_21(i*32 + 2) + x_30(i*32 + 3) + x_38(i*32 + 4) + x_46(i*32 + 5) + x_53(i*32 + 6) + x_60(i*32 + 7) + x_66(i*32 + 8) + x_72(i*32 + 9) + x_77(i*32 + 10) + x_80(i*32 + 11) + x_84(i*32 + 12) + x_86(i*32 + 13) + x_88(i*32 + 14) + x_90(i*32 + 15) + x_90(i*32 + 16) + x_89(i*32 + 17) + x_87(i*32 + 18) + x_85(i*32 + 19) + x_82(i*32 + 20) + x_78(i*32 + 21) + x_74(i*32 + 22) + x_68(i*32 + 23) + x_63(i*32 + 24) + x_56(i*32 + 25) + x_50(i*32 + 26) + x_42(i*32 + 27) + x_34(i*32 + 28) + x_26(i*32 + 29) + x_17(i*32 + 30) + x_9(i*32 + 31);
						y_dst(i*32 + 1) <= x_9(i*32 + 0) + x_26(i*32 + 1) + x_42(i*32 + 2) + x_56(i*32 + 3) + x_68(i*32 + 4) + x_78(i*32 + 5) + x_85(i*32 + 6) + x_89(i*32 + 7) + x_90(i*32 + 8) + x_86(i*32 + 9) + x_80(i*32 + 10) + x_72(i*32 + 11) + x_60(i*32 + 12) + x_46(i*32 + 13) + x_30(i*32 + 14) + x_13(i*32 + 15) - x_4(i*32 + 16) - x_21(i*32 + 17) - x_38(i*32 + 18) - x_53(i*32 + 19) - x_66(i*32 + 20) - x_77(i*32 + 21) - x_84(i*32 + 22) - x_88(i*32 + 23) - x_90(i*32 + 24) - x_87(i*32 + 25) - x_82(i*32 + 26) - x_74(i*32 + 27) - x_63(i*32 + 28) - x_50(i*32 + 29) - x_34(i*32 + 30) - x_17(i*32 + 31);
						y_dst(i*32 + 2) <= x_13(i*32 + 0) + x_38(i*32 + 1) + x_60(i*32 + 2) + x_77(i*32 + 3) + x_86(i*32 + 4) + x_90(i*32 + 5) + x_85(i*32 + 6) + x_74(i*32 + 7) + x_56(i*32 + 8) + x_34(i*32 + 9) + x_9(i*32 + 10) - x_17(i*32 + 11) - x_42(i*32 + 12) - x_63(i*32 + 13) - x_78(i*32 + 14) - x_87(i*32 + 15) - x_90(i*32 + 16) - x_84(i*32 + 17) - x_72(i*32 + 18) - x_53(i*32 + 19) - x_30(i*32 + 20) - x_4(i*32 + 21) + x_21(i*32 + 22) + x_46(i*32 + 23) + x_66(i*32 + 24) + x_80(i*32 + 25) + x_88(i*32 + 26) + x_89(i*32 + 27) + x_82(i*32 + 28) + x_68(i*32 + 29) + x_50(i*32 + 30) + x_26(i*32 + 31);
						y_dst(i*32 + 3) <= x_17(i*32 + 0) + x_50(i*32 + 1) + x_74(i*32 + 2) + x_87(i*32 + 3) + x_88(i*32 + 4) + x_77(i*32 + 5) + x_53(i*32 + 6) + x_21(i*32 + 7) - x_13(i*32 + 8) - x_46(i*32 + 9) - x_72(i*32 + 10) - x_86(i*32 + 11) - x_89(i*32 + 12) - x_78(i*32 + 13) - x_56(i*32 + 14) - x_26(i*32 + 15) + x_9(i*32 + 16) + x_42(i*32 + 17) + x_68(i*32 + 18) + x_85(i*32 + 19) + x_90(i*32 + 20) + x_80(i*32 + 21) + x_60(i*32 + 22) + x_30(i*32 + 23) - x_4(i*32 + 24) - x_38(i*32 + 25) - x_66(i*32 + 26) - x_84(i*32 + 27) - x_90(i*32 + 28) - x_82(i*32 + 29) - x_63(i*32 + 30) - x_34(i*32 + 31);
						y_dst(i*32 + 4) <= x_21(i*32 + 0) + x_60(i*32 + 1) + x_84(i*32 + 2) + x_89(i*32 + 3) + x_74(i*32 + 4) + x_42(i*32 + 5) - x_42(i*32 + 7) - x_74(i*32 + 8) - x_89(i*32 + 9) - x_84(i*32 + 10) - x_60(i*32 + 11) - x_21(i*32 + 12) + x_21(i*32 + 13) + x_60(i*32 + 14) + x_84(i*32 + 15) + x_89(i*32 + 16) + x_74(i*32 + 17) + x_42(i*32 + 18) - x_42(i*32 + 20) - x_74(i*32 + 21) - x_89(i*32 + 22) - x_84(i*32 + 23) - x_60(i*32 + 24) - x_21(i*32 + 25) + x_21(i*32 + 26) + x_60(i*32 + 27) + x_84(i*32 + 28) + x_89(i*32 + 29) + x_74(i*32 + 30) + x_42(i*32 + 31);
						y_dst(i*32 + 5) <= x_26(i*32 + 0) + x_68(i*32 + 1) + x_89(i*32 + 2) + x_80(i*32 + 3) + x_46(i*32 + 4) - x_4(i*32 + 5) - x_53(i*32 + 6) - x_84(i*32 + 7) - x_87(i*32 + 8) - x_63(i*32 + 9) - x_17(i*32 + 10) + x_34(i*32 + 11) + x_74(i*32 + 12) + x_90(i*32 + 13) + x_77(i*32 + 14) + x_38(i*32 + 15) - x_13(i*32 + 16) - x_60(i*32 + 17) - x_86(i*32 + 18) - x_85(i*32 + 19) - x_56(i*32 + 20) - x_9(i*32 + 21) + x_42(i*32 + 22) + x_78(i*32 + 23) + x_90(i*32 + 24) + x_72(i*32 + 25) + x_30(i*32 + 26) - x_21(i*32 + 27) - x_66(i*32 + 28) - x_88(i*32 + 29) - x_82(i*32 + 30) - x_50(i*32 + 31);
						y_dst(i*32 + 6) <= x_30(i*32 + 0) + x_77(i*32 + 1) + x_89(i*32 + 2) + x_63(i*32 + 3) + x_9(i*32 + 4) - x_50(i*32 + 5) - x_85(i*32 + 6) - x_84(i*32 + 7) - x_46(i*32 + 8) + x_13(i*32 + 9) + x_66(i*32 + 10) + x_90(i*32 + 11) + x_74(i*32 + 12) + x_26(i*32 + 13) - x_34(i*32 + 14) - x_78(i*32 + 15) - x_88(i*32 + 16) - x_60(i*32 + 17) - x_4(i*32 + 18) + x_53(i*32 + 19) + x_86(i*32 + 20) + x_82(i*32 + 21) + x_42(i*32 + 22) - x_17(i*32 + 23) - x_68(i*32 + 24) - x_90(i*32 + 25) - x_72(i*32 + 26) - x_21(i*32 + 27) + x_38(i*32 + 28) + x_80(i*32 + 29) + x_87(i*32 + 30) + x_56(i*32 + 31);
						y_dst(i*32 + 7) <= x_34(i*32 + 0) + x_82(i*32 + 1) + x_84(i*32 + 2) + x_38(i*32 + 3) - x_30(i*32 + 4) - x_80(i*32 + 5) - x_85(i*32 + 6) - x_42(i*32 + 7) + x_26(i*32 + 8) + x_78(i*32 + 9) + x_86(i*32 + 10) + x_46(i*32 + 11) - x_21(i*32 + 12) - x_77(i*32 + 13) - x_87(i*32 + 14) - x_50(i*32 + 15) + x_17(i*32 + 16) + x_74(i*32 + 17) + x_88(i*32 + 18) + x_53(i*32 + 19) - x_13(i*32 + 20) - x_72(i*32 + 21) - x_89(i*32 + 22) - x_56(i*32 + 23) + x_9(i*32 + 24) + x_68(i*32 + 25) + x_90(i*32 + 26) + x_60(i*32 + 27) - x_4(i*32 + 28) - x_66(i*32 + 29) - x_90(i*32 + 30) - x_63(i*32 + 31);
						y_dst(i*32 + 8) <= x_38(i*32 + 0) + x_86(i*32 + 1) + x_74(i*32 + 2) + x_9(i*32 + 3) - x_63(i*32 + 4) - x_90(i*32 + 5) - x_53(i*32 + 6) + x_21(i*32 + 7) + x_80(i*32 + 8) + x_82(i*32 + 9) + x_26(i*32 + 10) - x_50(i*32 + 11) - x_89(i*32 + 12) - x_66(i*32 + 13) + x_4(i*32 + 14) + x_72(i*32 + 15) + x_87(i*32 + 16) + x_42(i*32 + 17) - x_34(i*32 + 18) - x_85(i*32 + 19) - x_77(i*32 + 20) - x_13(i*32 + 21) + x_60(i*32 + 22) + x_90(i*32 + 23) + x_56(i*32 + 24) - x_17(i*32 + 25) - x_78(i*32 + 26) - x_84(i*32 + 27) - x_30(i*32 + 28) + x_46(i*32 + 29) + x_88(i*32 + 30) + x_68(i*32 + 31);
						y_dst(i*32 + 9) <= x_42(i*32 + 0) + x_89(i*32 + 1) + x_60(i*32 + 2) - x_21(i*32 + 3) - x_84(i*32 + 4) - x_74(i*32 + 5) + x_74(i*32 + 7) + x_84(i*32 + 8) + x_21(i*32 + 9) - x_60(i*32 + 10) - x_89(i*32 + 11) - x_42(i*32 + 12) + x_42(i*32 + 13) + x_89(i*32 + 14) + x_60(i*32 + 15) - x_21(i*32 + 16) - x_84(i*32 + 17) - x_74(i*32 + 18) + x_74(i*32 + 20) + x_84(i*32 + 21) + x_21(i*32 + 22) - x_60(i*32 + 23) - x_89(i*32 + 24) - x_42(i*32 + 25) + x_42(i*32 + 26) + x_89(i*32 + 27) + x_60(i*32 + 28) - x_21(i*32 + 29) - x_84(i*32 + 30) - x_74(i*32 + 31);
						y_dst(i*32 + 10) <= x_46(i*32 + 0) + x_90(i*32 + 1) + x_42(i*32 + 2) - x_50(i*32 + 3) - x_90(i*32 + 4) - x_38(i*32 + 5) + x_53(i*32 + 6) + x_89(i*32 + 7) + x_34(i*32 + 8) - x_56(i*32 + 9) - x_88(i*32 + 10) - x_30(i*32 + 11) + x_60(i*32 + 12) + x_87(i*32 + 13) + x_26(i*32 + 14) - x_63(i*32 + 15) - x_86(i*32 + 16) - x_21(i*32 + 17) + x_66(i*32 + 18) + x_85(i*32 + 19) + x_17(i*32 + 20) - x_68(i*32 + 21) - x_84(i*32 + 22) - x_13(i*32 + 23) + x_72(i*32 + 24) + x_82(i*32 + 25) + x_9(i*32 + 26) - x_74(i*32 + 27) - x_80(i*32 + 28) - x_4(i*32 + 29) + x_77(i*32 + 30) + x_78(i*32 + 31);
						y_dst(i*32 + 11) <= x_50(i*32 + 0) + x_88(i*32 + 1) + x_21(i*32 + 2) - x_72(i*32 + 3) - x_78(i*32 + 4) + x_9(i*32 + 5) + x_85(i*32 + 6) + x_60(i*32 + 7) - x_38(i*32 + 8) - x_90(i*32 + 9) - x_34(i*32 + 10) + x_63(i*32 + 11) + x_84(i*32 + 12) + x_4(i*32 + 13) - x_80(i*32 + 14) - x_68(i*32 + 15) + x_26(i*32 + 16) + x_89(i*32 + 17) + x_46(i*32 + 18) - x_53(i*32 + 19) - x_87(i*32 + 20) - x_17(i*32 + 21) + x_74(i*32 + 22) + x_77(i*32 + 23) - x_13(i*32 + 24) - x_86(i*32 + 25) - x_56(i*32 + 26) + x_42(i*32 + 27) + x_90(i*32 + 28) + x_30(i*32 + 29) - x_66(i*32 + 30) - x_82(i*32 + 31);
						y_dst(i*32 + 12) <= x_53(i*32 + 0) + x_85(i*32 + 1) - x_85(i*32 + 3) - x_53(i*32 + 4) + x_53(i*32 + 5) + x_85(i*32 + 6) - x_85(i*32 + 8) - x_53(i*32 + 9) + x_53(i*32 + 10) + x_85(i*32 + 11) - x_85(i*32 + 13) - x_53(i*32 + 14) + x_53(i*32 + 15) + x_85(i*32 + 16) - x_85(i*32 + 18) - x_53(i*32 + 19) + x_53(i*32 + 20) + x_85(i*32 + 21) - x_85(i*32 + 23) - x_53(i*32 + 24) + x_53(i*32 + 25) + x_85(i*32 + 26) - x_85(i*32 + 28) - x_53(i*32 + 29) + x_53(i*32 + 30) + x_85(i*32 + 31);
						y_dst(i*32 + 13) <= x_56(i*32 + 0) + x_80(i*32 + 1) - x_21(i*32 + 2) - x_90(i*32 + 3) - x_17(i*32 + 4) + x_82(i*32 + 5) + x_53(i*32 + 6) - x_60(i*32 + 7) - x_78(i*32 + 8) + x_26(i*32 + 9) + x_90(i*32 + 10) + x_13(i*32 + 11) - x_84(i*32 + 12) - x_50(i*32 + 13) + x_63(i*32 + 14) + x_77(i*32 + 15) - x_30(i*32 + 16) - x_89(i*32 + 17) - x_9(i*32 + 18) + x_85(i*32 + 19) + x_46(i*32 + 20) - x_66(i*32 + 21) - x_74(i*32 + 22) + x_34(i*32 + 23) + x_88(i*32 + 24) + x_4(i*32 + 25) - x_86(i*32 + 26) - x_42(i*32 + 27) + x_68(i*32 + 28) + x_72(i*32 + 29) - x_38(i*32 + 30) - x_87(i*32 + 31);
						y_dst(i*32 + 14) <= x_60(i*32 + 0) + x_74(i*32 + 1) - x_42(i*32 + 2) - x_84(i*32 + 3) + x_21(i*32 + 4) + x_89(i*32 + 5) - x_89(i*32 + 7) - x_21(i*32 + 8) + x_84(i*32 + 9) + x_42(i*32 + 10) - x_74(i*32 + 11) - x_60(i*32 + 12) + x_60(i*32 + 13) + x_74(i*32 + 14) - x_42(i*32 + 15) - x_84(i*32 + 16) + x_21(i*32 + 17) + x_89(i*32 + 18) - x_89(i*32 + 20) - x_21(i*32 + 21) + x_84(i*32 + 22) + x_42(i*32 + 23) - x_74(i*32 + 24) - x_60(i*32 + 25) + x_60(i*32 + 26) + x_74(i*32 + 27) - x_42(i*32 + 28) - x_84(i*32 + 29) + x_21(i*32 + 30) + x_89(i*32 + 31);
						y_dst(i*32 + 15) <= x_63(i*32 + 0) + x_66(i*32 + 1) - x_60(i*32 + 2) - x_68(i*32 + 3) + x_56(i*32 + 4) + x_72(i*32 + 5) - x_53(i*32 + 6) - x_74(i*32 + 7) + x_50(i*32 + 8) + x_77(i*32 + 9) - x_46(i*32 + 10) - x_78(i*32 + 11) + x_42(i*32 + 12) + x_80(i*32 + 13) - x_38(i*32 + 14) - x_82(i*32 + 15) + x_34(i*32 + 16) + x_84(i*32 + 17) - x_30(i*32 + 18) - x_85(i*32 + 19) + x_26(i*32 + 20) + x_86(i*32 + 21) - x_21(i*32 + 22) - x_87(i*32 + 23) + x_17(i*32 + 24) + x_88(i*32 + 25) - x_13(i*32 + 26) - x_89(i*32 + 27) + x_9(i*32 + 28) + x_90(i*32 + 29) - x_4(i*32 + 30) - x_90(i*32 + 31);
						y_dst(i*32 + 16) <= x_66(i*32 + 0) + x_56(i*32 + 1) - x_74(i*32 + 2) - x_46(i*32 + 3) + x_80(i*32 + 4) + x_34(i*32 + 5) - x_85(i*32 + 6) - x_21(i*32 + 7) + x_88(i*32 + 8) + x_9(i*32 + 9) - x_90(i*32 + 10) + x_4(i*32 + 11) + x_89(i*32 + 12) - x_17(i*32 + 13) - x_86(i*32 + 14) + x_30(i*32 + 15) + x_82(i*32 + 16) - x_42(i*32 + 17) - x_77(i*32 + 18) + x_53(i*32 + 19) + x_68(i*32 + 20) - x_63(i*32 + 21) - x_60(i*32 + 22) + x_72(i*32 + 23) + x_50(i*32 + 24) - x_78(i*32 + 25) - x_38(i*32 + 26) + x_84(i*32 + 27) + x_26(i*32 + 28) - x_87(i*32 + 29) - x_13(i*32 + 30) + x_90(i*32 + 31);
						y_dst(i*32 + 17) <= x_68(i*32 + 0) + x_46(i*32 + 1) - x_84(i*32 + 2) - x_17(i*32 + 3) + x_90(i*32 + 4) - x_13(i*32 + 5) - x_85(i*32 + 6) + x_42(i*32 + 7) + x_72(i*32 + 8) - x_66(i*32 + 9) - x_50(i*32 + 10) + x_82(i*32 + 11) + x_21(i*32 + 12) - x_90(i*32 + 13) + x_9(i*32 + 14) + x_86(i*32 + 15) - x_38(i*32 + 16) - x_74(i*32 + 17) + x_63(i*32 + 18) + x_53(i*32 + 19) - x_80(i*32 + 20) - x_26(i*32 + 21) + x_89(i*32 + 22) - x_4(i*32 + 23) - x_87(i*32 + 24) + x_34(i*32 + 25) + x_77(i*32 + 26) - x_60(i*32 + 27) - x_56(i*32 + 28) + x_78(i*32 + 29) + x_30(i*32 + 30) - x_88(i*32 + 31);
						y_dst(i*32 + 18) <= x_72(i*32 + 0) + x_34(i*32 + 1) - x_89(i*32 + 2) + x_13(i*32 + 3) + x_82(i*32 + 4) - x_56(i*32 + 5) - x_53(i*32 + 6) + x_84(i*32 + 7) + x_9(i*32 + 8) - x_88(i*32 + 9) + x_38(i*32 + 10) + x_68(i*32 + 11) - x_74(i*32 + 12) - x_30(i*32 + 13) + x_90(i*32 + 14) - x_17(i*32 + 15) - x_80(i*32 + 16) + x_60(i*32 + 17) + x_50(i*32 + 18) - x_85(i*32 + 19) - x_4(i*32 + 20) + x_87(i*32 + 21) - x_42(i*32 + 22) - x_66(i*32 + 23) + x_77(i*32 + 24) + x_26(i*32 + 25) - x_90(i*32 + 26) + x_21(i*32 + 27) + x_78(i*32 + 28) - x_63(i*32 + 29) - x_46(i*32 + 30) + x_86(i*32 + 31);
						y_dst(i*32 + 19) <= x_74(i*32 + 0) + x_21(i*32 + 1) - x_89(i*32 + 2) + x_42(i*32 + 3) + x_60(i*32 + 4) - x_84(i*32 + 5) + x_84(i*32 + 7) - x_60(i*32 + 8) - x_42(i*32 + 9) + x_89(i*32 + 10) - x_21(i*32 + 11) - x_74(i*32 + 12) + x_74(i*32 + 13) + x_21(i*32 + 14) - x_89(i*32 + 15) + x_42(i*32 + 16) + x_60(i*32 + 17) - x_84(i*32 + 18) + x_84(i*32 + 20) - x_60(i*32 + 21) - x_42(i*32 + 22) + x_89(i*32 + 23) - x_21(i*32 + 24) - x_74(i*32 + 25) + x_74(i*32 + 26) + x_21(i*32 + 27) - x_89(i*32 + 28) + x_42(i*32 + 29) + x_60(i*32 + 30) - x_84(i*32 + 31);
						y_dst(i*32 + 20) <= x_77(i*32 + 0) + x_9(i*32 + 1) - x_84(i*32 + 2) + x_66(i*32 + 3) + x_26(i*32 + 4) - x_88(i*32 + 5) + x_53(i*32 + 6) + x_42(i*32 + 7) - x_90(i*32 + 8) + x_38(i*32 + 9) + x_56(i*32 + 10) - x_87(i*32 + 11) + x_21(i*32 + 12) + x_68(i*32 + 13) - x_82(i*32 + 14) + x_4(i*32 + 15) + x_78(i*32 + 16) - x_74(i*32 + 17) - x_13(i*32 + 18) + x_85(i*32 + 19) - x_63(i*32 + 20) - x_30(i*32 + 21) + x_89(i*32 + 22) - x_50(i*32 + 23) - x_46(i*32 + 24) + x_90(i*32 + 25) - x_34(i*32 + 26) - x_60(i*32 + 27) + x_86(i*32 + 28) - x_17(i*32 + 29) - x_72(i*32 + 30) + x_80(i*32 + 31);
						y_dst(i*32 + 21) <= x_78(i*32 + 0) - x_4(i*32 + 1) - x_74(i*32 + 2) + x_82(i*32 + 3) - x_13(i*32 + 4) - x_68(i*32 + 5) + x_85(i*32 + 6) - x_21(i*32 + 7) - x_63(i*32 + 8) + x_87(i*32 + 9) - x_30(i*32 + 10) - x_56(i*32 + 11) + x_89(i*32 + 12) - x_38(i*32 + 13) - x_50(i*32 + 14) + x_90(i*32 + 15) - x_46(i*32 + 16) - x_42(i*32 + 17) + x_90(i*32 + 18) - x_53(i*32 + 19) - x_34(i*32 + 20) + x_88(i*32 + 21) - x_60(i*32 + 22) - x_26(i*32 + 23) + x_86(i*32 + 24) - x_66(i*32 + 25) - x_17(i*32 + 26) + x_84(i*32 + 27) - x_72(i*32 + 28) - x_9(i*32 + 29) + x_80(i*32 + 30) - x_77(i*32 + 31);
						y_dst(i*32 + 22) <= x_80(i*32 + 0) - x_17(i*32 + 1) - x_60(i*32 + 2) + x_90(i*32 + 3) - x_50(i*32 + 4) - x_30(i*32 + 5) + x_85(i*32 + 6) - x_74(i*32 + 7) + x_4(i*32 + 8) + x_68(i*32 + 9) - x_87(i*32 + 10) + x_38(i*32 + 11) + x_42(i*32 + 12) - x_88(i*32 + 13) + x_66(i*32 + 14) + x_9(i*32 + 15) - x_77(i*32 + 16) + x_84(i*32 + 17) - x_26(i*32 + 18) - x_53(i*32 + 19) + x_90(i*32 + 20) - x_56(i*32 + 21) - x_21(i*32 + 22) + x_82(i*32 + 23) - x_78(i*32 + 24) + x_13(i*32 + 25) + x_63(i*32 + 26) - x_89(i*32 + 27) + x_46(i*32 + 28) + x_34(i*32 + 29) - x_86(i*32 + 30) + x_72(i*32 + 31);
						y_dst(i*32 + 23) <= x_82(i*32 + 0) - x_30(i*32 + 1) - x_42(i*32 + 2) + x_86(i*32 + 3) - x_77(i*32 + 4) + x_17(i*32 + 5) + x_53(i*32 + 6) - x_89(i*32 + 7) + x_68(i*32 + 8) - x_4(i*32 + 9) - x_63(i*32 + 10) + x_90(i*32 + 11) - x_60(i*32 + 12) - x_9(i*32 + 13) + x_72(i*32 + 14) - x_88(i*32 + 15) + x_50(i*32 + 16) + x_21(i*32 + 17) - x_78(i*32 + 18) + x_85(i*32 + 19) - x_38(i*32 + 20) - x_34(i*32 + 21) + x_84(i*32 + 22) - x_80(i*32 + 23) + x_26(i*32 + 24) + x_46(i*32 + 25) - x_87(i*32 + 26) + x_74(i*32 + 27) - x_13(i*32 + 28) - x_56(i*32 + 29) + x_90(i*32 + 30) - x_66(i*32 + 31);
						y_dst(i*32 + 24) <= x_84(i*32 + 0) - x_42(i*32 + 1) - x_21(i*32 + 2) + x_74(i*32 + 3) - x_89(i*32 + 4) + x_60(i*32 + 5) - x_60(i*32 + 7) + x_89(i*32 + 8) - x_74(i*32 + 9) + x_21(i*32 + 10) + x_42(i*32 + 11) - x_84(i*32 + 12) + x_84(i*32 + 13) - x_42(i*32 + 14) - x_21(i*32 + 15) + x_74(i*32 + 16) - x_89(i*32 + 17) + x_60(i*32 + 18) - x_60(i*32 + 20) + x_89(i*32 + 21) - x_74(i*32 + 22) + x_21(i*32 + 23) + x_42(i*32 + 24) - x_84(i*32 + 25) + x_84(i*32 + 26) - x_42(i*32 + 27) - x_21(i*32 + 28) + x_74(i*32 + 29) - x_89(i*32 + 30) + x_60(i*32 + 31);
						y_dst(i*32 + 25) <= x_85(i*32 + 0) - x_53(i*32 + 1) + x_53(i*32 + 3) - x_85(i*32 + 4) + x_85(i*32 + 5) - x_53(i*32 + 6) + x_53(i*32 + 8) - x_85(i*32 + 9) + x_85(i*32 + 10) - x_53(i*32 + 11) + x_53(i*32 + 13) - x_85(i*32 + 14) + x_85(i*32 + 15) - x_53(i*32 + 16) + x_53(i*32 + 18) - x_85(i*32 + 19) + x_85(i*32 + 20) - x_53(i*32 + 21) + x_53(i*32 + 23) - x_85(i*32 + 24) + x_85(i*32 + 25) - x_53(i*32 + 26) + x_53(i*32 + 28) - x_85(i*32 + 29) + x_85(i*32 + 30) - x_53(i*32 + 31);
						y_dst(i*32 + 26) <= x_86(i*32 + 0) - x_63(i*32 + 1) + x_21(i*32 + 2) + x_26(i*32 + 3) - x_66(i*32 + 4) + x_87(i*32 + 5) - x_85(i*32 + 6) + x_60(i*32 + 7) - x_17(i*32 + 8) - x_30(i*32 + 9) + x_68(i*32 + 10) - x_88(i*32 + 11) + x_84(i*32 + 12) - x_56(i*32 + 13) + x_13(i*32 + 14) + x_34(i*32 + 15) - x_72(i*32 + 16) + x_89(i*32 + 17) - x_82(i*32 + 18) + x_53(i*32 + 19) - x_9(i*32 + 20) - x_38(i*32 + 21) + x_74(i*32 + 22) - x_90(i*32 + 23) + x_80(i*32 + 24) - x_50(i*32 + 25) + x_4(i*32 + 26) + x_42(i*32 + 27) - x_77(i*32 + 28) + x_90(i*32 + 29) - x_78(i*32 + 30) + x_46(i*32 + 31);
						y_dst(i*32 + 27) <= x_87(i*32 + 0) - x_72(i*32 + 1) + x_42(i*32 + 2) - x_4(i*32 + 3) - x_34(i*32 + 4) + x_66(i*32 + 5) - x_85(i*32 + 6) + x_89(i*32 + 7) - x_77(i*32 + 8) + x_50(i*32 + 9) - x_13(i*32 + 10) - x_26(i*32 + 11) + x_60(i*32 + 12) - x_82(i*32 + 13) + x_90(i*32 + 14) - x_80(i*32 + 15) + x_56(i*32 + 16) - x_21(i*32 + 17) - x_17(i*32 + 18) + x_53(i*32 + 19) - x_78(i*32 + 20) + x_90(i*32 + 21) - x_84(i*32 + 22) + x_63(i*32 + 23) - x_30(i*32 + 24) - x_9(i*32 + 25) + x_46(i*32 + 26) - x_74(i*32 + 27) + x_88(i*32 + 28) - x_86(i*32 + 29) + x_68(i*32 + 30) - x_38(i*32 + 31);
						y_dst(i*32 + 28) <= x_88(i*32 + 0) - x_78(i*32 + 1) + x_60(i*32 + 2) - x_34(i*32 + 3) + x_4(i*32 + 4) + x_26(i*32 + 5) - x_53(i*32 + 6) + x_74(i*32 + 7) - x_86(i*32 + 8) + x_90(i*32 + 9) - x_82(i*32 + 10) + x_66(i*32 + 11) - x_42(i*32 + 12) + x_13(i*32 + 13) + x_17(i*32 + 14) - x_46(i*32 + 15) + x_68(i*32 + 16) - x_84(i*32 + 17) + x_90(i*32 + 18) - x_85(i*32 + 19) + x_72(i*32 + 20) - x_50(i*32 + 21) + x_21(i*32 + 22) + x_9(i*32 + 23) - x_38(i*32 + 24) + x_63(i*32 + 25) - x_80(i*32 + 26) + x_89(i*32 + 27) - x_87(i*32 + 28) + x_77(i*32 + 29) - x_56(i*32 + 30) + x_30(i*32 + 31);
						y_dst(i*32 + 29) <= x_89(i*32 + 0) - x_84(i*32 + 1) + x_74(i*32 + 2) - x_60(i*32 + 3) + x_42(i*32 + 4) - x_21(i*32 + 5) + x_21(i*32 + 7) - x_42(i*32 + 8) + x_60(i*32 + 9) - x_74(i*32 + 10) + x_84(i*32 + 11) - x_89(i*32 + 12) + x_89(i*32 + 13) - x_84(i*32 + 14) + x_74(i*32 + 15) - x_60(i*32 + 16) + x_42(i*32 + 17) - x_21(i*32 + 18) + x_21(i*32 + 20) - x_42(i*32 + 21) + x_60(i*32 + 22) - x_74(i*32 + 23) + x_84(i*32 + 24) - x_89(i*32 + 25) + x_89(i*32 + 26) - x_84(i*32 + 27) + x_74(i*32 + 28) - x_60(i*32 + 29) + x_42(i*32 + 30) - x_21(i*32 + 31);
						y_dst(i*32 + 30) <= x_90(i*32 + 0) - x_87(i*32 + 1) + x_84(i*32 + 2) - x_78(i*32 + 3) + x_72(i*32 + 4) - x_63(i*32 + 5) + x_53(i*32 + 6) - x_42(i*32 + 7) + x_30(i*32 + 8) - x_17(i*32 + 9) + x_4(i*32 + 10) + x_9(i*32 + 11) - x_21(i*32 + 12) + x_34(i*32 + 13) - x_46(i*32 + 14) + x_56(i*32 + 15) - x_66(i*32 + 16) + x_74(i*32 + 17) - x_80(i*32 + 18) + x_85(i*32 + 19) - x_88(i*32 + 20) + x_90(i*32 + 21) - x_89(i*32 + 22) + x_86(i*32 + 23) - x_82(i*32 + 24) + x_77(i*32 + 25) - x_68(i*32 + 26) + x_60(i*32 + 27) - x_50(i*32 + 28) + x_38(i*32 + 29) - x_26(i*32 + 30) + x_13(i*32 + 31);
						y_dst(i*32 + 31) <= x_90(i*32 + 0) - x_90(i*32 + 1) + x_89(i*32 + 2) - x_88(i*32 + 3) + x_87(i*32 + 4) - x_86(i*32 + 5) + x_85(i*32 + 6) - x_84(i*32 + 7) + x_82(i*32 + 8) - x_80(i*32 + 9) + x_78(i*32 + 10) - x_77(i*32 + 11) + x_74(i*32 + 12) - x_72(i*32 + 13) + x_68(i*32 + 14) - x_66(i*32 + 15) + x_63(i*32 + 16) - x_60(i*32 + 17) + x_56(i*32 + 18) - x_53(i*32 + 19) + x_50(i*32 + 20) - x_46(i*32 + 21) + x_42(i*32 + 22) - x_38(i*32 + 23) + x_34(i*32 + 24) - x_30(i*32 + 25) + x_26(i*32 + 26) - x_21(i*32 + 27) + x_17(i*32 + 28) - x_13(i*32 + 29) + x_9(i*32 + 30) - x_4(i*32 + 31);
 
            end generate generateSignalsOutputsDST7;
				
			with op select
			y <= y_dct when '0',
			     y_dst when others;
        
y0 <= y(0);
y1 <= y(1);
y2 <= y(2);
y3 <= y(3);
y4 <= y(4);
y5 <= y(5);
y6 <= y(6);
y7 <= y(7);
y8 <= y(8);
y9 <= y(9);
y10 <= y(10);
y11 <= y(11);
y12 <= y(12);
y13 <= y(13);
y14 <= y(14);
y15 <= y(15);
y16 <= y(16);
y17 <= y(17);
y18 <= y(18);
y19 <= y(19);
y20 <= y(20);
y21 <= y(21);
y22 <= y(22);
y23 <= y(23);
y24 <= y(24);
y25 <= y(25);
y26 <= y(26);
y27 <= y(27);
y28 <= y(28);
y29 <= y(29);
y30 <= y(30);
y31 <= y(31);
y32 <= y(32);
y33 <= y(33);
y34 <= y(34);
y35 <= y(35);
y36 <= y(36);
y37 <= y(37);
y38 <= y(38);
y39 <= y(39);
y40 <= y(40);
y41 <= y(41);
y42 <= y(42);
y43 <= y(43);
y44 <= y(44);
y45 <= y(45);
y46 <= y(46);
y47 <= y(47);
y48 <= y(48);
y49 <= y(49);
y50 <= y(50);
y51 <= y(51);
y52 <= y(52);
y53 <= y(53);
y54 <= y(54);
y55 <= y(55);
y56 <= y(56);
y57 <= y(57);
y58 <= y(58);
y59 <= y(59);
y60 <= y(60);
y61 <= y(61);
y62 <= y(62);
y63 <= y(63);
			

			
end behavior;
